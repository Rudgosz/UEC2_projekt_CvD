module game_fsm (
    input  logic clk,
    input  logic rst,
    input  logic enter_pressed_local,
    input  logic enter_pressed_remote,
    input  logic turn_done,
    input  logic [9:0] hp_local,
    input  logic [9:0] hp_remote,
    output logic whose_turn,
	output logic [2:0] state_game_fsm
);

    typedef enum logic [2:0] {
        START_SCREEN   = 3'b000,
        PLAYER_TURN    = 3'b001,
        OPPONENT_TURN  = 3'b010,
        CHECK_WIN      = 3'b011,
		GAME_OVER      = 3'b100
	} state_t;
	state_t state;

	assign state_game_fsm = state;

	always_ff @(posedge clk) begin
		if (rst) begin
			state       <= START_SCREEN;
			whose_turn  <= 0;
		end else begin
			case (state)

				START_SCREEN: begin
					if (enter_pressed_local) begin
						whose_turn <= 1;
						state <= PLAYER_TURN;
					end else if (enter_pressed_remote) begin
						whose_turn <= 0;
						state <= OPPONENT_TURN;
					end
				end

				PLAYER_TURN: begin
					whose_turn <= 1;
					if (turn_done) begin
						whose_turn <= 0;
						state <= CHECK_WIN;
					end
				end

				OPPONENT_TURN: begin
					whose_turn <= 0;
					if (turn_done) begin
						whose_turn <= 1;
						state <= CHECK_WIN;
					end
				end

				CHECK_WIN: begin
					if (hp_local == 0 || hp_remote == 0) begin
						state <= GAME_OVER;
					end else if (whose_turn) begin
						whose_turn <= 1;
						state <= PLAYER_TURN;
					end else begin
						whose_turn <= 0;
						state <= OPPONENT_TURN;
					end
				end

				GAME_OVER: begin
					whose_turn <= 0; // no one's turn
					if (enter_pressed_local || enter_pressed_remote)
						state <= START_SCREEN;
				end

				default: begin
					state <= START_SCREEN;
					whose_turn <= 0;
				end
			endcase
		end
	end


endmodule